module mod(a, d);

input wire [324:0] a;
output wire [164:0] d;

assign d[0:7]       = a[0:7]    ^a[163:170] ^a[317:324] ^a[279:286] ^a[246:253];                                                                            //5
assign d[8]         = a[8]      ^a[171]     ^a[287]     ^a[254];                                                                                            //4
assign d[9:16]      = a[9:16]   ^a[172:179] ^a[163:170] ^a[317:324] ^a[288:295] ^a[279:286] ^a[255:262] ^a[246:253];                                        //8
assign d[17:45]     = a[17:45]  ^a[180:208] ^a[171:199] ^a[296:324] ^a[287:315] ^a[263:291] ^a[254:282];                                                    //7
assign d[46]        = a[46]     ^a[209]     ^a[200]     ^a[316]     ^a[292]     ^a[283];                                                                    //6
assign d[47:54]     = a[47:54]  ^a[210:217] ^a[201:208] ^a[163:170] ^a[317:324] ^a[317:324] ^a[279:286] ^a[293:300] ^a[284:291] ^a[246:253];                //10
assign d[55:78]     = a[55:78]  ^a[218:241] ^a[209:232] ^a[171:194] ^a[287:310] ^a[301:324] ^a[292:315] ^a[254:277];                                        //8
assign d[79]        = a[79]     ^a[242]     ^a[233]     ^a[195]     ^a[311]     ^a[316]     ^a[278];                                                        //7
assign d[80:87]     = a[80:87]  ^a[243:250] ^a[234:241] ^a[196:203] ^a[163:170] ^a[317:324] ^a[312:319] ^a[279:286] ^a[317:324] ^a[279:286] ^a[246:253];    //11
assign d[88:92]     = a[88:92]  ^a[251:255] ^a[242:246] ^a[204:208] ^a[171:175] ^a[320:324] ^a[287:291] ^a[287:291] ^a[254:258];                            //9
assign d[93:125]    = a[93:125] ^a[256:288] ^a[247:279] ^a[209:241] ^a[176:208] ^a[292:324] ^a[292:324] ^a[259:291];                                        //8
assign d[126:158]   = a[126:158]^a[289:321] ^a[280:312] ^a[242:274] ^a[209:241] ^a[292:324];                                                                //6
assign d[159:161]   = a[159:161]^a[322:324] ^a[313:315] ^a[275:277] ^a[242:244];                                                                            //5
assign d[162]       = a[162]    ^a[316]     ^a[278]     ^a[245];                                                                                            //4

endmodule